// nios_security.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module nios_security (
		input  wire        clk_clk,        //     clk.clk
		output wire [31:0] duty_export,    //    duty.export
		output wire [31:0] led0_export,    //    led0.export
		output wire        led1_export,    //    led1.export
		output wire        led2_export,    //    led2.export
		output wire        led3_export,    //    led3.export
		output wire        led4_export,    //    led4.export
		output wire        led5_export,    //    led5.export
		output wire        led6_export,    //    led6.export
		output wire        led7_export,    //    led7.export
		output wire        led8_export,    //    led8.export
		output wire        led9_export,    //    led9.export
		output wire [31:0] period_export,  //  period.export
		input  wire        pwm_in_export,  //  pwm_in.export
		output wire        pwm_out_export, // pwm_out.export
		input  wire        reset_reset_n,  //   reset.reset_n
		output wire [31:0] stop_export,    //    stop.export
		input  wire        sw_export,      //      sw.export
		input  wire        uart_rxd,       //    uart.rxd
		output wire        uart_txd        //        .txd
	);

	wire  [31:0] niosii_data_master_readdata;                          // mm_interconnect_0:NIOSII_data_master_readdata -> NIOSII:d_readdata
	wire         niosii_data_master_waitrequest;                       // mm_interconnect_0:NIOSII_data_master_waitrequest -> NIOSII:d_waitrequest
	wire         niosii_data_master_debugaccess;                       // NIOSII:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:NIOSII_data_master_debugaccess
	wire  [18:0] niosii_data_master_address;                           // NIOSII:d_address -> mm_interconnect_0:NIOSII_data_master_address
	wire   [3:0] niosii_data_master_byteenable;                        // NIOSII:d_byteenable -> mm_interconnect_0:NIOSII_data_master_byteenable
	wire         niosii_data_master_read;                              // NIOSII:d_read -> mm_interconnect_0:NIOSII_data_master_read
	wire         niosii_data_master_write;                             // NIOSII:d_write -> mm_interconnect_0:NIOSII_data_master_write
	wire  [31:0] niosii_data_master_writedata;                         // NIOSII:d_writedata -> mm_interconnect_0:NIOSII_data_master_writedata
	wire  [31:0] niosii_instruction_master_readdata;                   // mm_interconnect_0:NIOSII_instruction_master_readdata -> NIOSII:i_readdata
	wire         niosii_instruction_master_waitrequest;                // mm_interconnect_0:NIOSII_instruction_master_waitrequest -> NIOSII:i_waitrequest
	wire  [18:0] niosii_instruction_master_address;                    // NIOSII:i_address -> mm_interconnect_0:NIOSII_instruction_master_address
	wire         niosii_instruction_master_read;                       // NIOSII:i_read -> mm_interconnect_0:NIOSII_instruction_master_read
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_chipselect;  // mm_interconnect_0:JTAG_avalon_jtag_slave_chipselect -> JTAG:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_readdata;    // JTAG:av_readdata -> mm_interconnect_0:JTAG_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest; // JTAG:av_waitrequest -> mm_interconnect_0:JTAG_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_avalon_jtag_slave_address;     // mm_interconnect_0:JTAG_avalon_jtag_slave_address -> JTAG:av_address
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_read;        // mm_interconnect_0:JTAG_avalon_jtag_slave_read -> JTAG:av_read_n
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_write;       // mm_interconnect_0:JTAG_avalon_jtag_slave_write -> JTAG:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_writedata;   // mm_interconnect_0:JTAG_avalon_jtag_slave_writedata -> JTAG:av_writedata
	wire  [31:0] mm_interconnect_0_id_control_slave_readdata;          // ID:readdata -> mm_interconnect_0:ID_control_slave_readdata
	wire   [0:0] mm_interconnect_0_id_control_slave_address;           // mm_interconnect_0:ID_control_slave_address -> ID:address
	wire  [31:0] mm_interconnect_0_niosii_debug_mem_slave_readdata;    // NIOSII:debug_mem_slave_readdata -> mm_interconnect_0:NIOSII_debug_mem_slave_readdata
	wire         mm_interconnect_0_niosii_debug_mem_slave_waitrequest; // NIOSII:debug_mem_slave_waitrequest -> mm_interconnect_0:NIOSII_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_niosii_debug_mem_slave_debugaccess; // mm_interconnect_0:NIOSII_debug_mem_slave_debugaccess -> NIOSII:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_niosii_debug_mem_slave_address;     // mm_interconnect_0:NIOSII_debug_mem_slave_address -> NIOSII:debug_mem_slave_address
	wire         mm_interconnect_0_niosii_debug_mem_slave_read;        // mm_interconnect_0:NIOSII_debug_mem_slave_read -> NIOSII:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_niosii_debug_mem_slave_byteenable;  // mm_interconnect_0:NIOSII_debug_mem_slave_byteenable -> NIOSII:debug_mem_slave_byteenable
	wire         mm_interconnect_0_niosii_debug_mem_slave_write;       // mm_interconnect_0:NIOSII_debug_mem_slave_write -> NIOSII:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_niosii_debug_mem_slave_writedata;   // mm_interconnect_0:NIOSII_debug_mem_slave_writedata -> NIOSII:debug_mem_slave_writedata
	wire         mm_interconnect_0_uart_s1_chipselect;                 // mm_interconnect_0:UART_s1_chipselect -> UART:chipselect
	wire  [15:0] mm_interconnect_0_uart_s1_readdata;                   // UART:readdata -> mm_interconnect_0:UART_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_s1_address;                    // mm_interconnect_0:UART_s1_address -> UART:address
	wire         mm_interconnect_0_uart_s1_read;                       // mm_interconnect_0:UART_s1_read -> UART:read_n
	wire         mm_interconnect_0_uart_s1_begintransfer;              // mm_interconnect_0:UART_s1_begintransfer -> UART:begintransfer
	wire         mm_interconnect_0_uart_s1_write;                      // mm_interconnect_0:UART_s1_write -> UART:write_n
	wire  [15:0] mm_interconnect_0_uart_s1_writedata;                  // mm_interconnect_0:UART_s1_writedata -> UART:writedata
	wire         mm_interconnect_0_ram_s1_chipselect;                  // mm_interconnect_0:RAM_s1_chipselect -> RAM:chipselect
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;                    // RAM:readdata -> mm_interconnect_0:RAM_s1_readdata
	wire  [14:0] mm_interconnect_0_ram_s1_address;                     // mm_interconnect_0:RAM_s1_address -> RAM:address
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;                  // mm_interconnect_0:RAM_s1_byteenable -> RAM:byteenable
	wire         mm_interconnect_0_ram_s1_write;                       // mm_interconnect_0:RAM_s1_write -> RAM:write
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;                   // mm_interconnect_0:RAM_s1_writedata -> RAM:writedata
	wire         mm_interconnect_0_ram_s1_clken;                       // mm_interconnect_0:RAM_s1_clken -> RAM:clken
	wire         mm_interconnect_0_stop_s1_chipselect;                 // mm_interconnect_0:STOP_s1_chipselect -> STOP:chipselect
	wire  [31:0] mm_interconnect_0_stop_s1_readdata;                   // STOP:readdata -> mm_interconnect_0:STOP_s1_readdata
	wire   [1:0] mm_interconnect_0_stop_s1_address;                    // mm_interconnect_0:STOP_s1_address -> STOP:address
	wire         mm_interconnect_0_stop_s1_write;                      // mm_interconnect_0:STOP_s1_write -> STOP:write_n
	wire  [31:0] mm_interconnect_0_stop_s1_writedata;                  // mm_interconnect_0:STOP_s1_writedata -> STOP:writedata
	wire         mm_interconnect_0_led0_s1_chipselect;                 // mm_interconnect_0:LED0_s1_chipselect -> LED0:chipselect
	wire  [31:0] mm_interconnect_0_led0_s1_readdata;                   // LED0:readdata -> mm_interconnect_0:LED0_s1_readdata
	wire   [1:0] mm_interconnect_0_led0_s1_address;                    // mm_interconnect_0:LED0_s1_address -> LED0:address
	wire         mm_interconnect_0_led0_s1_write;                      // mm_interconnect_0:LED0_s1_write -> LED0:write_n
	wire  [31:0] mm_interconnect_0_led0_s1_writedata;                  // mm_interconnect_0:LED0_s1_writedata -> LED0:writedata
	wire         mm_interconnect_0_duty_s1_chipselect;                 // mm_interconnect_0:DUTY_s1_chipselect -> DUTY:chipselect
	wire  [31:0] mm_interconnect_0_duty_s1_readdata;                   // DUTY:readdata -> mm_interconnect_0:DUTY_s1_readdata
	wire   [1:0] mm_interconnect_0_duty_s1_address;                    // mm_interconnect_0:DUTY_s1_address -> DUTY:address
	wire         mm_interconnect_0_duty_s1_write;                      // mm_interconnect_0:DUTY_s1_write -> DUTY:write_n
	wire  [31:0] mm_interconnect_0_duty_s1_writedata;                  // mm_interconnect_0:DUTY_s1_writedata -> DUTY:writedata
	wire         mm_interconnect_0_period_s1_chipselect;               // mm_interconnect_0:PERIOD_s1_chipselect -> PERIOD:chipselect
	wire  [31:0] mm_interconnect_0_period_s1_readdata;                 // PERIOD:readdata -> mm_interconnect_0:PERIOD_s1_readdata
	wire   [1:0] mm_interconnect_0_period_s1_address;                  // mm_interconnect_0:PERIOD_s1_address -> PERIOD:address
	wire         mm_interconnect_0_period_s1_write;                    // mm_interconnect_0:PERIOD_s1_write -> PERIOD:write_n
	wire  [31:0] mm_interconnect_0_period_s1_writedata;                // mm_interconnect_0:PERIOD_s1_writedata -> PERIOD:writedata
	wire  [31:0] mm_interconnect_0_sw_s1_readdata;                     // SW:readdata -> mm_interconnect_0:SW_s1_readdata
	wire   [1:0] mm_interconnect_0_sw_s1_address;                      // mm_interconnect_0:SW_s1_address -> SW:address
	wire  [31:0] mm_interconnect_0_pwm_in_s1_readdata;                 // PWM_IN:readdata -> mm_interconnect_0:PWM_IN_s1_readdata
	wire   [1:0] mm_interconnect_0_pwm_in_s1_address;                  // mm_interconnect_0:PWM_IN_s1_address -> PWM_IN:address
	wire         mm_interconnect_0_pwm_out_s1_chipselect;              // mm_interconnect_0:PWM_OUT_s1_chipselect -> PWM_OUT:chipselect
	wire  [31:0] mm_interconnect_0_pwm_out_s1_readdata;                // PWM_OUT:readdata -> mm_interconnect_0:PWM_OUT_s1_readdata
	wire   [1:0] mm_interconnect_0_pwm_out_s1_address;                 // mm_interconnect_0:PWM_OUT_s1_address -> PWM_OUT:address
	wire         mm_interconnect_0_pwm_out_s1_write;                   // mm_interconnect_0:PWM_OUT_s1_write -> PWM_OUT:write_n
	wire  [31:0] mm_interconnect_0_pwm_out_s1_writedata;               // mm_interconnect_0:PWM_OUT_s1_writedata -> PWM_OUT:writedata
	wire         mm_interconnect_0_led1_s1_chipselect;                 // mm_interconnect_0:LED1_s1_chipselect -> LED1:chipselect
	wire  [31:0] mm_interconnect_0_led1_s1_readdata;                   // LED1:readdata -> mm_interconnect_0:LED1_s1_readdata
	wire   [1:0] mm_interconnect_0_led1_s1_address;                    // mm_interconnect_0:LED1_s1_address -> LED1:address
	wire         mm_interconnect_0_led1_s1_write;                      // mm_interconnect_0:LED1_s1_write -> LED1:write_n
	wire  [31:0] mm_interconnect_0_led1_s1_writedata;                  // mm_interconnect_0:LED1_s1_writedata -> LED1:writedata
	wire         mm_interconnect_0_led7_s1_chipselect;                 // mm_interconnect_0:LED7_s1_chipselect -> LED7:chipselect
	wire  [31:0] mm_interconnect_0_led7_s1_readdata;                   // LED7:readdata -> mm_interconnect_0:LED7_s1_readdata
	wire   [1:0] mm_interconnect_0_led7_s1_address;                    // mm_interconnect_0:LED7_s1_address -> LED7:address
	wire         mm_interconnect_0_led7_s1_write;                      // mm_interconnect_0:LED7_s1_write -> LED7:write_n
	wire  [31:0] mm_interconnect_0_led7_s1_writedata;                  // mm_interconnect_0:LED7_s1_writedata -> LED7:writedata
	wire         mm_interconnect_0_led6_s1_chipselect;                 // mm_interconnect_0:LED6_s1_chipselect -> LED6:chipselect
	wire  [31:0] mm_interconnect_0_led6_s1_readdata;                   // LED6:readdata -> mm_interconnect_0:LED6_s1_readdata
	wire   [1:0] mm_interconnect_0_led6_s1_address;                    // mm_interconnect_0:LED6_s1_address -> LED6:address
	wire         mm_interconnect_0_led6_s1_write;                      // mm_interconnect_0:LED6_s1_write -> LED6:write_n
	wire  [31:0] mm_interconnect_0_led6_s1_writedata;                  // mm_interconnect_0:LED6_s1_writedata -> LED6:writedata
	wire         mm_interconnect_0_led5_s1_chipselect;                 // mm_interconnect_0:LED5_s1_chipselect -> LED5:chipselect
	wire  [31:0] mm_interconnect_0_led5_s1_readdata;                   // LED5:readdata -> mm_interconnect_0:LED5_s1_readdata
	wire   [1:0] mm_interconnect_0_led5_s1_address;                    // mm_interconnect_0:LED5_s1_address -> LED5:address
	wire         mm_interconnect_0_led5_s1_write;                      // mm_interconnect_0:LED5_s1_write -> LED5:write_n
	wire  [31:0] mm_interconnect_0_led5_s1_writedata;                  // mm_interconnect_0:LED5_s1_writedata -> LED5:writedata
	wire         mm_interconnect_0_led4_s1_chipselect;                 // mm_interconnect_0:LED4_s1_chipselect -> LED4:chipselect
	wire  [31:0] mm_interconnect_0_led4_s1_readdata;                   // LED4:readdata -> mm_interconnect_0:LED4_s1_readdata
	wire   [1:0] mm_interconnect_0_led4_s1_address;                    // mm_interconnect_0:LED4_s1_address -> LED4:address
	wire         mm_interconnect_0_led4_s1_write;                      // mm_interconnect_0:LED4_s1_write -> LED4:write_n
	wire  [31:0] mm_interconnect_0_led4_s1_writedata;                  // mm_interconnect_0:LED4_s1_writedata -> LED4:writedata
	wire         mm_interconnect_0_led3_s1_chipselect;                 // mm_interconnect_0:LED3_s1_chipselect -> LED3:chipselect
	wire  [31:0] mm_interconnect_0_led3_s1_readdata;                   // LED3:readdata -> mm_interconnect_0:LED3_s1_readdata
	wire   [1:0] mm_interconnect_0_led3_s1_address;                    // mm_interconnect_0:LED3_s1_address -> LED3:address
	wire         mm_interconnect_0_led3_s1_write;                      // mm_interconnect_0:LED3_s1_write -> LED3:write_n
	wire  [31:0] mm_interconnect_0_led3_s1_writedata;                  // mm_interconnect_0:LED3_s1_writedata -> LED3:writedata
	wire         mm_interconnect_0_led2_s1_chipselect;                 // mm_interconnect_0:LED2_s1_chipselect -> LED2:chipselect
	wire  [31:0] mm_interconnect_0_led2_s1_readdata;                   // LED2:readdata -> mm_interconnect_0:LED2_s1_readdata
	wire   [1:0] mm_interconnect_0_led2_s1_address;                    // mm_interconnect_0:LED2_s1_address -> LED2:address
	wire         mm_interconnect_0_led2_s1_write;                      // mm_interconnect_0:LED2_s1_write -> LED2:write_n
	wire  [31:0] mm_interconnect_0_led2_s1_writedata;                  // mm_interconnect_0:LED2_s1_writedata -> LED2:writedata
	wire         mm_interconnect_0_led8_s1_chipselect;                 // mm_interconnect_0:LED8_s1_chipselect -> LED8:chipselect
	wire  [31:0] mm_interconnect_0_led8_s1_readdata;                   // LED8:readdata -> mm_interconnect_0:LED8_s1_readdata
	wire   [1:0] mm_interconnect_0_led8_s1_address;                    // mm_interconnect_0:LED8_s1_address -> LED8:address
	wire         mm_interconnect_0_led8_s1_write;                      // mm_interconnect_0:LED8_s1_write -> LED8:write_n
	wire  [31:0] mm_interconnect_0_led8_s1_writedata;                  // mm_interconnect_0:LED8_s1_writedata -> LED8:writedata
	wire         mm_interconnect_0_led9_s1_chipselect;                 // mm_interconnect_0:LED9_s1_chipselect -> LED9:chipselect
	wire  [31:0] mm_interconnect_0_led9_s1_readdata;                   // LED9:readdata -> mm_interconnect_0:LED9_s1_readdata
	wire   [1:0] mm_interconnect_0_led9_s1_address;                    // mm_interconnect_0:LED9_s1_address -> LED9:address
	wire         mm_interconnect_0_led9_s1_write;                      // mm_interconnect_0:LED9_s1_write -> LED9:write_n
	wire  [31:0] mm_interconnect_0_led9_s1_writedata;                  // mm_interconnect_0:LED9_s1_writedata -> LED9:writedata
	wire         irq_mapper_receiver0_irq;                             // UART:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                             // JTAG:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] niosii_irq_irq;                                       // irq_mapper:sender_irq -> NIOSII:irq
	wire         rst_controller_reset_out_reset;                       // rst_controller:reset_out -> [DUTY:reset_n, ID:reset_n, JTAG:rst_n, LED0:reset_n, LED1:reset_n, LED2:reset_n, LED3:reset_n, LED4:reset_n, LED5:reset_n, LED6:reset_n, LED7:reset_n, LED8:reset_n, LED9:reset_n, NIOSII:reset_n, PERIOD:reset_n, PWM_IN:reset_n, PWM_OUT:reset_n, RAM:reset, STOP:reset_n, SW:reset_n, UART:reset_n, irq_mapper:reset, mm_interconnect_0:NIOSII_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                   // rst_controller:reset_req -> [NIOSII:reset_req, RAM:reset_req, rst_translator:reset_req_in]
	wire         niosii_debug_reset_request_reset;                     // NIOSII:debug_reset_request -> rst_controller:reset_in1

	nios_security_DUTY duty (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_duty_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_duty_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_duty_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_duty_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_duty_s1_readdata),   //                    .readdata
		.out_port   (duty_export)                           // external_connection.export
	);

	nios_security_ID id (
		.clock    (clk_clk),                                     //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),             //         reset.reset_n
		.readdata (mm_interconnect_0_id_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_id_control_slave_address)   //              .address
	);

	nios_security_JTAG jtag (
		.clk            (clk_clk),                                              //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                      //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                              //               irq.irq
	);

	nios_security_DUTY led0 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_led0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led0_s1_readdata),   //                    .readdata
		.out_port   (led0_export)                           // external_connection.export
	);

	nios_security_LED1 led1 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_led1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led1_s1_readdata),   //                    .readdata
		.out_port   (led1_export)                           // external_connection.export
	);

	nios_security_LED1 led2 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_led2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led2_s1_readdata),   //                    .readdata
		.out_port   (led2_export)                           // external_connection.export
	);

	nios_security_LED1 led3 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_led3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led3_s1_readdata),   //                    .readdata
		.out_port   (led3_export)                           // external_connection.export
	);

	nios_security_LED1 led4 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_led4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led4_s1_readdata),   //                    .readdata
		.out_port   (led4_export)                           // external_connection.export
	);

	nios_security_LED1 led5 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_led5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led5_s1_readdata),   //                    .readdata
		.out_port   (led5_export)                           // external_connection.export
	);

	nios_security_LED1 led6 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_led6_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led6_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led6_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led6_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led6_s1_readdata),   //                    .readdata
		.out_port   (led6_export)                           // external_connection.export
	);

	nios_security_LED1 led7 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_led7_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led7_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led7_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led7_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led7_s1_readdata),   //                    .readdata
		.out_port   (led7_export)                           // external_connection.export
	);

	nios_security_LED1 led8 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_led8_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led8_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led8_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led8_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led8_s1_readdata),   //                    .readdata
		.out_port   (led8_export)                           // external_connection.export
	);

	nios_security_LED1 led9 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_led9_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led9_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led9_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led9_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led9_s1_readdata),   //                    .readdata
		.out_port   (led9_export)                           // external_connection.export
	);

	nios_security_NIOSII niosii (
		.clk                                 (clk_clk),                                              //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                      //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                   //                          .reset_req
		.d_address                           (niosii_data_master_address),                           //               data_master.address
		.d_byteenable                        (niosii_data_master_byteenable),                        //                          .byteenable
		.d_read                              (niosii_data_master_read),                              //                          .read
		.d_readdata                          (niosii_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (niosii_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (niosii_data_master_write),                             //                          .write
		.d_writedata                         (niosii_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (niosii_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (niosii_instruction_master_address),                    //        instruction_master.address
		.i_read                              (niosii_instruction_master_read),                       //                          .read
		.i_readdata                          (niosii_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (niosii_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (niosii_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (niosii_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_niosii_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_niosii_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_niosii_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_niosii_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_niosii_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_niosii_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_niosii_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_niosii_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                      // custom_instruction_master.readra
	);

	nios_security_DUTY period (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_period_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_period_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_period_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_period_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_period_s1_readdata),   //                    .readdata
		.out_port   (period_export)                           // external_connection.export
	);

	nios_security_PWM_IN pwm_in (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_pwm_in_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pwm_in_s1_readdata), //                    .readdata
		.in_port  (pwm_in_export)                         // external_connection.export
	);

	nios_security_LED1 pwm_out (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_pwm_out_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pwm_out_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pwm_out_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pwm_out_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pwm_out_s1_readdata),   //                    .readdata
		.out_port   (pwm_out_export)                           // external_connection.export
	);

	nios_security_RAM ram (
		.clk        (clk_clk),                             //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze     (1'b0)                                 // (terminated)
	);

	nios_security_DUTY stop (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_stop_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_stop_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_stop_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_stop_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_stop_s1_readdata),   //                    .readdata
		.out_port   (stop_export)                           // external_connection.export
	);

	nios_security_PWM_IN sw (
		.clk      (clk_clk),                          //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),  //               reset.reset_n
		.address  (mm_interconnect_0_sw_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sw_s1_readdata), //                    .readdata
		.in_port  (sw_export)                         // external_connection.export
	);

	nios_security_UART uart (
		.clk           (clk_clk),                                 //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address       (mm_interconnect_0_uart_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_s1_readdata),      //                    .readdata
		.rxd           (uart_rxd),                                // external_connection.export
		.txd           (uart_txd),                                //                    .export
		.irq           (irq_mapper_receiver0_irq)                 //                 irq.irq
	);

	nios_security_mm_interconnect_0 mm_interconnect_0 (
		.CLK_clk_clk                              (clk_clk),                                              //                            CLK_clk.clk
		.NIOSII_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                       // NIOSII_reset_reset_bridge_in_reset.reset
		.NIOSII_data_master_address               (niosii_data_master_address),                           //                 NIOSII_data_master.address
		.NIOSII_data_master_waitrequest           (niosii_data_master_waitrequest),                       //                                   .waitrequest
		.NIOSII_data_master_byteenable            (niosii_data_master_byteenable),                        //                                   .byteenable
		.NIOSII_data_master_read                  (niosii_data_master_read),                              //                                   .read
		.NIOSII_data_master_readdata              (niosii_data_master_readdata),                          //                                   .readdata
		.NIOSII_data_master_write                 (niosii_data_master_write),                             //                                   .write
		.NIOSII_data_master_writedata             (niosii_data_master_writedata),                         //                                   .writedata
		.NIOSII_data_master_debugaccess           (niosii_data_master_debugaccess),                       //                                   .debugaccess
		.NIOSII_instruction_master_address        (niosii_instruction_master_address),                    //          NIOSII_instruction_master.address
		.NIOSII_instruction_master_waitrequest    (niosii_instruction_master_waitrequest),                //                                   .waitrequest
		.NIOSII_instruction_master_read           (niosii_instruction_master_read),                       //                                   .read
		.NIOSII_instruction_master_readdata       (niosii_instruction_master_readdata),                   //                                   .readdata
		.DUTY_s1_address                          (mm_interconnect_0_duty_s1_address),                    //                            DUTY_s1.address
		.DUTY_s1_write                            (mm_interconnect_0_duty_s1_write),                      //                                   .write
		.DUTY_s1_readdata                         (mm_interconnect_0_duty_s1_readdata),                   //                                   .readdata
		.DUTY_s1_writedata                        (mm_interconnect_0_duty_s1_writedata),                  //                                   .writedata
		.DUTY_s1_chipselect                       (mm_interconnect_0_duty_s1_chipselect),                 //                                   .chipselect
		.ID_control_slave_address                 (mm_interconnect_0_id_control_slave_address),           //                   ID_control_slave.address
		.ID_control_slave_readdata                (mm_interconnect_0_id_control_slave_readdata),          //                                   .readdata
		.JTAG_avalon_jtag_slave_address           (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //             JTAG_avalon_jtag_slave.address
		.JTAG_avalon_jtag_slave_write             (mm_interconnect_0_jtag_avalon_jtag_slave_write),       //                                   .write
		.JTAG_avalon_jtag_slave_read              (mm_interconnect_0_jtag_avalon_jtag_slave_read),        //                                   .read
		.JTAG_avalon_jtag_slave_readdata          (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                                   .readdata
		.JTAG_avalon_jtag_slave_writedata         (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                                   .writedata
		.JTAG_avalon_jtag_slave_waitrequest       (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                                   .waitrequest
		.JTAG_avalon_jtag_slave_chipselect        (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  //                                   .chipselect
		.LED0_s1_address                          (mm_interconnect_0_led0_s1_address),                    //                            LED0_s1.address
		.LED0_s1_write                            (mm_interconnect_0_led0_s1_write),                      //                                   .write
		.LED0_s1_readdata                         (mm_interconnect_0_led0_s1_readdata),                   //                                   .readdata
		.LED0_s1_writedata                        (mm_interconnect_0_led0_s1_writedata),                  //                                   .writedata
		.LED0_s1_chipselect                       (mm_interconnect_0_led0_s1_chipselect),                 //                                   .chipselect
		.LED1_s1_address                          (mm_interconnect_0_led1_s1_address),                    //                            LED1_s1.address
		.LED1_s1_write                            (mm_interconnect_0_led1_s1_write),                      //                                   .write
		.LED1_s1_readdata                         (mm_interconnect_0_led1_s1_readdata),                   //                                   .readdata
		.LED1_s1_writedata                        (mm_interconnect_0_led1_s1_writedata),                  //                                   .writedata
		.LED1_s1_chipselect                       (mm_interconnect_0_led1_s1_chipselect),                 //                                   .chipselect
		.LED2_s1_address                          (mm_interconnect_0_led2_s1_address),                    //                            LED2_s1.address
		.LED2_s1_write                            (mm_interconnect_0_led2_s1_write),                      //                                   .write
		.LED2_s1_readdata                         (mm_interconnect_0_led2_s1_readdata),                   //                                   .readdata
		.LED2_s1_writedata                        (mm_interconnect_0_led2_s1_writedata),                  //                                   .writedata
		.LED2_s1_chipselect                       (mm_interconnect_0_led2_s1_chipselect),                 //                                   .chipselect
		.LED3_s1_address                          (mm_interconnect_0_led3_s1_address),                    //                            LED3_s1.address
		.LED3_s1_write                            (mm_interconnect_0_led3_s1_write),                      //                                   .write
		.LED3_s1_readdata                         (mm_interconnect_0_led3_s1_readdata),                   //                                   .readdata
		.LED3_s1_writedata                        (mm_interconnect_0_led3_s1_writedata),                  //                                   .writedata
		.LED3_s1_chipselect                       (mm_interconnect_0_led3_s1_chipselect),                 //                                   .chipselect
		.LED4_s1_address                          (mm_interconnect_0_led4_s1_address),                    //                            LED4_s1.address
		.LED4_s1_write                            (mm_interconnect_0_led4_s1_write),                      //                                   .write
		.LED4_s1_readdata                         (mm_interconnect_0_led4_s1_readdata),                   //                                   .readdata
		.LED4_s1_writedata                        (mm_interconnect_0_led4_s1_writedata),                  //                                   .writedata
		.LED4_s1_chipselect                       (mm_interconnect_0_led4_s1_chipselect),                 //                                   .chipselect
		.LED5_s1_address                          (mm_interconnect_0_led5_s1_address),                    //                            LED5_s1.address
		.LED5_s1_write                            (mm_interconnect_0_led5_s1_write),                      //                                   .write
		.LED5_s1_readdata                         (mm_interconnect_0_led5_s1_readdata),                   //                                   .readdata
		.LED5_s1_writedata                        (mm_interconnect_0_led5_s1_writedata),                  //                                   .writedata
		.LED5_s1_chipselect                       (mm_interconnect_0_led5_s1_chipselect),                 //                                   .chipselect
		.LED6_s1_address                          (mm_interconnect_0_led6_s1_address),                    //                            LED6_s1.address
		.LED6_s1_write                            (mm_interconnect_0_led6_s1_write),                      //                                   .write
		.LED6_s1_readdata                         (mm_interconnect_0_led6_s1_readdata),                   //                                   .readdata
		.LED6_s1_writedata                        (mm_interconnect_0_led6_s1_writedata),                  //                                   .writedata
		.LED6_s1_chipselect                       (mm_interconnect_0_led6_s1_chipselect),                 //                                   .chipselect
		.LED7_s1_address                          (mm_interconnect_0_led7_s1_address),                    //                            LED7_s1.address
		.LED7_s1_write                            (mm_interconnect_0_led7_s1_write),                      //                                   .write
		.LED7_s1_readdata                         (mm_interconnect_0_led7_s1_readdata),                   //                                   .readdata
		.LED7_s1_writedata                        (mm_interconnect_0_led7_s1_writedata),                  //                                   .writedata
		.LED7_s1_chipselect                       (mm_interconnect_0_led7_s1_chipselect),                 //                                   .chipselect
		.LED8_s1_address                          (mm_interconnect_0_led8_s1_address),                    //                            LED8_s1.address
		.LED8_s1_write                            (mm_interconnect_0_led8_s1_write),                      //                                   .write
		.LED8_s1_readdata                         (mm_interconnect_0_led8_s1_readdata),                   //                                   .readdata
		.LED8_s1_writedata                        (mm_interconnect_0_led8_s1_writedata),                  //                                   .writedata
		.LED8_s1_chipselect                       (mm_interconnect_0_led8_s1_chipselect),                 //                                   .chipselect
		.LED9_s1_address                          (mm_interconnect_0_led9_s1_address),                    //                            LED9_s1.address
		.LED9_s1_write                            (mm_interconnect_0_led9_s1_write),                      //                                   .write
		.LED9_s1_readdata                         (mm_interconnect_0_led9_s1_readdata),                   //                                   .readdata
		.LED9_s1_writedata                        (mm_interconnect_0_led9_s1_writedata),                  //                                   .writedata
		.LED9_s1_chipselect                       (mm_interconnect_0_led9_s1_chipselect),                 //                                   .chipselect
		.NIOSII_debug_mem_slave_address           (mm_interconnect_0_niosii_debug_mem_slave_address),     //             NIOSII_debug_mem_slave.address
		.NIOSII_debug_mem_slave_write             (mm_interconnect_0_niosii_debug_mem_slave_write),       //                                   .write
		.NIOSII_debug_mem_slave_read              (mm_interconnect_0_niosii_debug_mem_slave_read),        //                                   .read
		.NIOSII_debug_mem_slave_readdata          (mm_interconnect_0_niosii_debug_mem_slave_readdata),    //                                   .readdata
		.NIOSII_debug_mem_slave_writedata         (mm_interconnect_0_niosii_debug_mem_slave_writedata),   //                                   .writedata
		.NIOSII_debug_mem_slave_byteenable        (mm_interconnect_0_niosii_debug_mem_slave_byteenable),  //                                   .byteenable
		.NIOSII_debug_mem_slave_waitrequest       (mm_interconnect_0_niosii_debug_mem_slave_waitrequest), //                                   .waitrequest
		.NIOSII_debug_mem_slave_debugaccess       (mm_interconnect_0_niosii_debug_mem_slave_debugaccess), //                                   .debugaccess
		.PERIOD_s1_address                        (mm_interconnect_0_period_s1_address),                  //                          PERIOD_s1.address
		.PERIOD_s1_write                          (mm_interconnect_0_period_s1_write),                    //                                   .write
		.PERIOD_s1_readdata                       (mm_interconnect_0_period_s1_readdata),                 //                                   .readdata
		.PERIOD_s1_writedata                      (mm_interconnect_0_period_s1_writedata),                //                                   .writedata
		.PERIOD_s1_chipselect                     (mm_interconnect_0_period_s1_chipselect),               //                                   .chipselect
		.PWM_IN_s1_address                        (mm_interconnect_0_pwm_in_s1_address),                  //                          PWM_IN_s1.address
		.PWM_IN_s1_readdata                       (mm_interconnect_0_pwm_in_s1_readdata),                 //                                   .readdata
		.PWM_OUT_s1_address                       (mm_interconnect_0_pwm_out_s1_address),                 //                         PWM_OUT_s1.address
		.PWM_OUT_s1_write                         (mm_interconnect_0_pwm_out_s1_write),                   //                                   .write
		.PWM_OUT_s1_readdata                      (mm_interconnect_0_pwm_out_s1_readdata),                //                                   .readdata
		.PWM_OUT_s1_writedata                     (mm_interconnect_0_pwm_out_s1_writedata),               //                                   .writedata
		.PWM_OUT_s1_chipselect                    (mm_interconnect_0_pwm_out_s1_chipselect),              //                                   .chipselect
		.RAM_s1_address                           (mm_interconnect_0_ram_s1_address),                     //                             RAM_s1.address
		.RAM_s1_write                             (mm_interconnect_0_ram_s1_write),                       //                                   .write
		.RAM_s1_readdata                          (mm_interconnect_0_ram_s1_readdata),                    //                                   .readdata
		.RAM_s1_writedata                         (mm_interconnect_0_ram_s1_writedata),                   //                                   .writedata
		.RAM_s1_byteenable                        (mm_interconnect_0_ram_s1_byteenable),                  //                                   .byteenable
		.RAM_s1_chipselect                        (mm_interconnect_0_ram_s1_chipselect),                  //                                   .chipselect
		.RAM_s1_clken                             (mm_interconnect_0_ram_s1_clken),                       //                                   .clken
		.STOP_s1_address                          (mm_interconnect_0_stop_s1_address),                    //                            STOP_s1.address
		.STOP_s1_write                            (mm_interconnect_0_stop_s1_write),                      //                                   .write
		.STOP_s1_readdata                         (mm_interconnect_0_stop_s1_readdata),                   //                                   .readdata
		.STOP_s1_writedata                        (mm_interconnect_0_stop_s1_writedata),                  //                                   .writedata
		.STOP_s1_chipselect                       (mm_interconnect_0_stop_s1_chipselect),                 //                                   .chipselect
		.SW_s1_address                            (mm_interconnect_0_sw_s1_address),                      //                              SW_s1.address
		.SW_s1_readdata                           (mm_interconnect_0_sw_s1_readdata),                     //                                   .readdata
		.UART_s1_address                          (mm_interconnect_0_uart_s1_address),                    //                            UART_s1.address
		.UART_s1_write                            (mm_interconnect_0_uart_s1_write),                      //                                   .write
		.UART_s1_read                             (mm_interconnect_0_uart_s1_read),                       //                                   .read
		.UART_s1_readdata                         (mm_interconnect_0_uart_s1_readdata),                   //                                   .readdata
		.UART_s1_writedata                        (mm_interconnect_0_uart_s1_writedata),                  //                                   .writedata
		.UART_s1_begintransfer                    (mm_interconnect_0_uart_s1_begintransfer),              //                                   .begintransfer
		.UART_s1_chipselect                       (mm_interconnect_0_uart_s1_chipselect)                  //                                   .chipselect
	);

	nios_security_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (niosii_irq_irq)                  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (niosii_debug_reset_request_reset),   // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule

// nios2e.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module nios2e (
		input  wire        clk_clk,       //   clk.clk
		output wire [27:0] cycle_export,  // cycle.export
		input  wire        dip0_export,   //  dip0.export
		input  wire [15:0] dip1_export,   //  dip1.export
		input  wire        dip2_export,   //  dip2.export
		input  wire        dip3_export,   //  dip3.export
		output wire [31:0] duty_export,   //  duty.export
		output wire        led0_export,   //  led0.export
		output wire        led1_export,   //  led1.export
		output wire        led2_export,   //  led2.export
		output wire        led3_export,   //  led3.export
		output wire        led4_export,   //  led4.export
		output wire        led5_export,   //  led5.export
		output wire        led6_export,   //  led6.export
		output wire        led7_export,   //  led7.export
		input  wire        reset_reset_n, // reset.reset_n
		input  wire [15:0] sw0_export,    //   sw0.export
		input  wire [15:0] sw1_export     //   sw1.export
	);

	wire  [31:0] nios2_data_master_readdata;                           // mm_interconnect_0:NIOS2_data_master_readdata -> NIOS2:d_readdata
	wire         nios2_data_master_waitrequest;                        // mm_interconnect_0:NIOS2_data_master_waitrequest -> NIOS2:d_waitrequest
	wire         nios2_data_master_debugaccess;                        // NIOS2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:NIOS2_data_master_debugaccess
	wire  [15:0] nios2_data_master_address;                            // NIOS2:d_address -> mm_interconnect_0:NIOS2_data_master_address
	wire   [3:0] nios2_data_master_byteenable;                         // NIOS2:d_byteenable -> mm_interconnect_0:NIOS2_data_master_byteenable
	wire         nios2_data_master_read;                               // NIOS2:d_read -> mm_interconnect_0:NIOS2_data_master_read
	wire         nios2_data_master_write;                              // NIOS2:d_write -> mm_interconnect_0:NIOS2_data_master_write
	wire  [31:0] nios2_data_master_writedata;                          // NIOS2:d_writedata -> mm_interconnect_0:NIOS2_data_master_writedata
	wire  [31:0] nios2_instruction_master_readdata;                    // mm_interconnect_0:NIOS2_instruction_master_readdata -> NIOS2:i_readdata
	wire         nios2_instruction_master_waitrequest;                 // mm_interconnect_0:NIOS2_instruction_master_waitrequest -> NIOS2:i_waitrequest
	wire  [15:0] nios2_instruction_master_address;                     // NIOS2:i_address -> mm_interconnect_0:NIOS2_instruction_master_address
	wire         nios2_instruction_master_read;                        // NIOS2:i_read -> mm_interconnect_0:NIOS2_instruction_master_read
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_chipselect;  // mm_interconnect_0:JTAG_avalon_jtag_slave_chipselect -> JTAG:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_readdata;    // JTAG:av_readdata -> mm_interconnect_0:JTAG_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest; // JTAG:av_waitrequest -> mm_interconnect_0:JTAG_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_avalon_jtag_slave_address;     // mm_interconnect_0:JTAG_avalon_jtag_slave_address -> JTAG:av_address
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_read;        // mm_interconnect_0:JTAG_avalon_jtag_slave_read -> JTAG:av_read_n
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_write;       // mm_interconnect_0:JTAG_avalon_jtag_slave_write -> JTAG:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_writedata;   // mm_interconnect_0:JTAG_avalon_jtag_slave_writedata -> JTAG:av_writedata
	wire  [31:0] mm_interconnect_0_id_control_slave_readdata;          // ID:readdata -> mm_interconnect_0:ID_control_slave_readdata
	wire   [0:0] mm_interconnect_0_id_control_slave_address;           // mm_interconnect_0:ID_control_slave_address -> ID:address
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_readdata;     // NIOS2:debug_mem_slave_readdata -> mm_interconnect_0:NIOS2_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_debug_mem_slave_waitrequest;  // NIOS2:debug_mem_slave_waitrequest -> mm_interconnect_0:NIOS2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_debug_mem_slave_debugaccess;  // mm_interconnect_0:NIOS2_debug_mem_slave_debugaccess -> NIOS2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_debug_mem_slave_address;      // mm_interconnect_0:NIOS2_debug_mem_slave_address -> NIOS2:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_debug_mem_slave_read;         // mm_interconnect_0:NIOS2_debug_mem_slave_read -> NIOS2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_debug_mem_slave_byteenable;   // mm_interconnect_0:NIOS2_debug_mem_slave_byteenable -> NIOS2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_debug_mem_slave_write;        // mm_interconnect_0:NIOS2_debug_mem_slave_write -> NIOS2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_writedata;    // mm_interconnect_0:NIOS2_debug_mem_slave_writedata -> NIOS2:debug_mem_slave_writedata
	wire         mm_interconnect_0_ram_s1_chipselect;                  // mm_interconnect_0:RAM_s1_chipselect -> RAM:chipselect
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;                    // RAM:readdata -> mm_interconnect_0:RAM_s1_readdata
	wire  [11:0] mm_interconnect_0_ram_s1_address;                     // mm_interconnect_0:RAM_s1_address -> RAM:address
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;                  // mm_interconnect_0:RAM_s1_byteenable -> RAM:byteenable
	wire         mm_interconnect_0_ram_s1_write;                       // mm_interconnect_0:RAM_s1_write -> RAM:write
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;                   // mm_interconnect_0:RAM_s1_writedata -> RAM:writedata
	wire         mm_interconnect_0_ram_s1_clken;                       // mm_interconnect_0:RAM_s1_clken -> RAM:clken
	wire         mm_interconnect_0_cycle_s1_chipselect;                // mm_interconnect_0:CYCLE_s1_chipselect -> CYCLE:chipselect
	wire  [31:0] mm_interconnect_0_cycle_s1_readdata;                  // CYCLE:readdata -> mm_interconnect_0:CYCLE_s1_readdata
	wire   [1:0] mm_interconnect_0_cycle_s1_address;                   // mm_interconnect_0:CYCLE_s1_address -> CYCLE:address
	wire         mm_interconnect_0_cycle_s1_write;                     // mm_interconnect_0:CYCLE_s1_write -> CYCLE:write_n
	wire  [31:0] mm_interconnect_0_cycle_s1_writedata;                 // mm_interconnect_0:CYCLE_s1_writedata -> CYCLE:writedata
	wire         mm_interconnect_0_duty_s1_chipselect;                 // mm_interconnect_0:DUTY_s1_chipselect -> DUTY:chipselect
	wire  [31:0] mm_interconnect_0_duty_s1_readdata;                   // DUTY:readdata -> mm_interconnect_0:DUTY_s1_readdata
	wire   [1:0] mm_interconnect_0_duty_s1_address;                    // mm_interconnect_0:DUTY_s1_address -> DUTY:address
	wire         mm_interconnect_0_duty_s1_write;                      // mm_interconnect_0:DUTY_s1_write -> DUTY:write_n
	wire  [31:0] mm_interconnect_0_duty_s1_writedata;                  // mm_interconnect_0:DUTY_s1_writedata -> DUTY:writedata
	wire  [31:0] mm_interconnect_0_dip1_s1_readdata;                   // DIP1:readdata -> mm_interconnect_0:DIP1_s1_readdata
	wire   [1:0] mm_interconnect_0_dip1_s1_address;                    // mm_interconnect_0:DIP1_s1_address -> DIP1:address
	wire  [31:0] mm_interconnect_0_sw1_s1_readdata;                    // SW1:readdata -> mm_interconnect_0:SW1_s1_readdata
	wire   [1:0] mm_interconnect_0_sw1_s1_address;                     // mm_interconnect_0:SW1_s1_address -> SW1:address
	wire  [31:0] mm_interconnect_0_sw0_s1_readdata;                    // SW0:readdata -> mm_interconnect_0:SW0_s1_readdata
	wire   [1:0] mm_interconnect_0_sw0_s1_address;                     // mm_interconnect_0:SW0_s1_address -> SW0:address
	wire         mm_interconnect_0_led1_s1_chipselect;                 // mm_interconnect_0:LED1_s1_chipselect -> LED1:chipselect
	wire  [31:0] mm_interconnect_0_led1_s1_readdata;                   // LED1:readdata -> mm_interconnect_0:LED1_s1_readdata
	wire   [1:0] mm_interconnect_0_led1_s1_address;                    // mm_interconnect_0:LED1_s1_address -> LED1:address
	wire         mm_interconnect_0_led1_s1_write;                      // mm_interconnect_0:LED1_s1_write -> LED1:write_n
	wire  [31:0] mm_interconnect_0_led1_s1_writedata;                  // mm_interconnect_0:LED1_s1_writedata -> LED1:writedata
	wire         mm_interconnect_0_led2_s1_chipselect;                 // mm_interconnect_0:LED2_s1_chipselect -> LED2:chipselect
	wire  [31:0] mm_interconnect_0_led2_s1_readdata;                   // LED2:readdata -> mm_interconnect_0:LED2_s1_readdata
	wire   [1:0] mm_interconnect_0_led2_s1_address;                    // mm_interconnect_0:LED2_s1_address -> LED2:address
	wire         mm_interconnect_0_led2_s1_write;                      // mm_interconnect_0:LED2_s1_write -> LED2:write_n
	wire  [31:0] mm_interconnect_0_led2_s1_writedata;                  // mm_interconnect_0:LED2_s1_writedata -> LED2:writedata
	wire         mm_interconnect_0_led3_s1_chipselect;                 // mm_interconnect_0:LED3_s1_chipselect -> LED3:chipselect
	wire  [31:0] mm_interconnect_0_led3_s1_readdata;                   // LED3:readdata -> mm_interconnect_0:LED3_s1_readdata
	wire   [1:0] mm_interconnect_0_led3_s1_address;                    // mm_interconnect_0:LED3_s1_address -> LED3:address
	wire         mm_interconnect_0_led3_s1_write;                      // mm_interconnect_0:LED3_s1_write -> LED3:write_n
	wire  [31:0] mm_interconnect_0_led3_s1_writedata;                  // mm_interconnect_0:LED3_s1_writedata -> LED3:writedata
	wire         mm_interconnect_0_led0_s1_chipselect;                 // mm_interconnect_0:LED0_s1_chipselect -> LED0:chipselect
	wire  [31:0] mm_interconnect_0_led0_s1_readdata;                   // LED0:readdata -> mm_interconnect_0:LED0_s1_readdata
	wire   [1:0] mm_interconnect_0_led0_s1_address;                    // mm_interconnect_0:LED0_s1_address -> LED0:address
	wire         mm_interconnect_0_led0_s1_write;                      // mm_interconnect_0:LED0_s1_write -> LED0:write_n
	wire  [31:0] mm_interconnect_0_led0_s1_writedata;                  // mm_interconnect_0:LED0_s1_writedata -> LED0:writedata
	wire  [31:0] mm_interconnect_0_dip3_s1_readdata;                   // DIP3:readdata -> mm_interconnect_0:DIP3_s1_readdata
	wire   [1:0] mm_interconnect_0_dip3_s1_address;                    // mm_interconnect_0:DIP3_s1_address -> DIP3:address
	wire  [31:0] mm_interconnect_0_dip2_s1_readdata;                   // DIP2:readdata -> mm_interconnect_0:DIP2_s1_readdata
	wire   [1:0] mm_interconnect_0_dip2_s1_address;                    // mm_interconnect_0:DIP2_s1_address -> DIP2:address
	wire  [31:0] mm_interconnect_0_dip0_s1_readdata;                   // DIP0:readdata -> mm_interconnect_0:DIP0_s1_readdata
	wire   [1:0] mm_interconnect_0_dip0_s1_address;                    // mm_interconnect_0:DIP0_s1_address -> DIP0:address
	wire         mm_interconnect_0_led4_s1_chipselect;                 // mm_interconnect_0:LED4_s1_chipselect -> LED4:chipselect
	wire  [31:0] mm_interconnect_0_led4_s1_readdata;                   // LED4:readdata -> mm_interconnect_0:LED4_s1_readdata
	wire   [1:0] mm_interconnect_0_led4_s1_address;                    // mm_interconnect_0:LED4_s1_address -> LED4:address
	wire         mm_interconnect_0_led4_s1_write;                      // mm_interconnect_0:LED4_s1_write -> LED4:write_n
	wire  [31:0] mm_interconnect_0_led4_s1_writedata;                  // mm_interconnect_0:LED4_s1_writedata -> LED4:writedata
	wire         mm_interconnect_0_led5_s1_chipselect;                 // mm_interconnect_0:LED5_s1_chipselect -> LED5:chipselect
	wire  [31:0] mm_interconnect_0_led5_s1_readdata;                   // LED5:readdata -> mm_interconnect_0:LED5_s1_readdata
	wire   [1:0] mm_interconnect_0_led5_s1_address;                    // mm_interconnect_0:LED5_s1_address -> LED5:address
	wire         mm_interconnect_0_led5_s1_write;                      // mm_interconnect_0:LED5_s1_write -> LED5:write_n
	wire  [31:0] mm_interconnect_0_led5_s1_writedata;                  // mm_interconnect_0:LED5_s1_writedata -> LED5:writedata
	wire         mm_interconnect_0_led7_s1_chipselect;                 // mm_interconnect_0:LED7_s1_chipselect -> LED7:chipselect
	wire  [31:0] mm_interconnect_0_led7_s1_readdata;                   // LED7:readdata -> mm_interconnect_0:LED7_s1_readdata
	wire   [1:0] mm_interconnect_0_led7_s1_address;                    // mm_interconnect_0:LED7_s1_address -> LED7:address
	wire         mm_interconnect_0_led7_s1_write;                      // mm_interconnect_0:LED7_s1_write -> LED7:write_n
	wire  [31:0] mm_interconnect_0_led7_s1_writedata;                  // mm_interconnect_0:LED7_s1_writedata -> LED7:writedata
	wire         mm_interconnect_0_led6_s1_chipselect;                 // mm_interconnect_0:LED6_s1_chipselect -> LED6:chipselect
	wire  [31:0] mm_interconnect_0_led6_s1_readdata;                   // LED6:readdata -> mm_interconnect_0:LED6_s1_readdata
	wire   [1:0] mm_interconnect_0_led6_s1_address;                    // mm_interconnect_0:LED6_s1_address -> LED6:address
	wire         mm_interconnect_0_led6_s1_write;                      // mm_interconnect_0:LED6_s1_write -> LED6:write_n
	wire  [31:0] mm_interconnect_0_led6_s1_writedata;                  // mm_interconnect_0:LED6_s1_writedata -> LED6:writedata
	wire         irq_mapper_receiver0_irq;                             // JTAG:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_irq_irq;                                        // irq_mapper:sender_irq -> NIOS2:irq
	wire         rst_controller_reset_out_reset;                       // rst_controller:reset_out -> [CYCLE:reset_n, DIP0:reset_n, DIP1:reset_n, DIP2:reset_n, DIP3:reset_n, DUTY:reset_n, ID:reset_n, JTAG:rst_n, LED0:reset_n, LED1:reset_n, LED2:reset_n, LED3:reset_n, LED4:reset_n, LED5:reset_n, LED6:reset_n, LED7:reset_n, NIOS2:reset_n, RAM:reset, SW0:reset_n, SW1:reset_n, irq_mapper:reset, mm_interconnect_0:NIOS2_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                   // rst_controller:reset_req -> [NIOS2:reset_req, RAM:reset_req, rst_translator:reset_req_in]
	wire         nios2_debug_reset_request_reset;                      // NIOS2:debug_reset_request -> rst_controller:reset_in1

	nios2e_CYCLE cycle (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_cycle_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_cycle_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_cycle_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_cycle_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_cycle_s1_readdata),   //                    .readdata
		.out_port   (cycle_export)                           // external_connection.export
	);

	nios2e_DIP0 dip0 (
		.clk      (clk_clk),                            //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address  (mm_interconnect_0_dip0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_dip0_s1_readdata), //                    .readdata
		.in_port  (dip0_export)                         // external_connection.export
	);

	nios2e_DIP1 dip1 (
		.clk      (clk_clk),                            //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address  (mm_interconnect_0_dip1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_dip1_s1_readdata), //                    .readdata
		.in_port  (dip1_export)                         // external_connection.export
	);

	nios2e_DIP0 dip2 (
		.clk      (clk_clk),                            //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address  (mm_interconnect_0_dip2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_dip2_s1_readdata), //                    .readdata
		.in_port  (dip2_export)                         // external_connection.export
	);

	nios2e_DIP0 dip3 (
		.clk      (clk_clk),                            //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address  (mm_interconnect_0_dip3_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_dip3_s1_readdata), //                    .readdata
		.in_port  (dip3_export)                         // external_connection.export
	);

	nios2e_DUTY duty (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_duty_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_duty_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_duty_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_duty_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_duty_s1_readdata),   //                    .readdata
		.out_port   (duty_export)                           // external_connection.export
	);

	nios2e_ID id (
		.clock    (clk_clk),                                     //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),             //         reset.reset_n
		.readdata (mm_interconnect_0_id_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_id_control_slave_address)   //              .address
	);

	nios2e_JTAG jtag (
		.clk            (clk_clk),                                              //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                      //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                              //               irq.irq
	);

	nios2e_LED0 led0 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_led0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led0_s1_readdata),   //                    .readdata
		.out_port   (led0_export)                           // external_connection.export
	);

	nios2e_LED0 led1 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_led1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led1_s1_readdata),   //                    .readdata
		.out_port   (led1_export)                           // external_connection.export
	);

	nios2e_LED0 led2 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_led2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led2_s1_readdata),   //                    .readdata
		.out_port   (led2_export)                           // external_connection.export
	);

	nios2e_LED0 led3 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_led3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led3_s1_readdata),   //                    .readdata
		.out_port   (led3_export)                           // external_connection.export
	);

	nios2e_LED0 led4 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_led4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led4_s1_readdata),   //                    .readdata
		.out_port   (led4_export)                           // external_connection.export
	);

	nios2e_LED0 led5 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_led5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led5_s1_readdata),   //                    .readdata
		.out_port   (led5_export)                           // external_connection.export
	);

	nios2e_LED0 led6 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_led6_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led6_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led6_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led6_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led6_s1_readdata),   //                    .readdata
		.out_port   (led6_export)                           // external_connection.export
	);

	nios2e_LED0 led7 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_led7_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led7_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led7_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led7_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led7_s1_readdata),   //                    .readdata
		.out_port   (led7_export)                           // external_connection.export
	);

	nios2e_NIOS2 nios2 (
		.clk                                 (clk_clk),                                             //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                     //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                           (nios2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_data_master_read),                              //                          .read
		.d_readdata                          (nios2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_data_master_write),                             //                          .write
		.d_writedata                         (nios2_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                     // custom_instruction_master.readra
	);

	nios2e_RAM ram (
		.clk        (clk_clk),                             //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze     (1'b0)                                 // (terminated)
	);

	nios2e_DIP1 sw0 (
		.clk      (clk_clk),                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),   //               reset.reset_n
		.address  (mm_interconnect_0_sw0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sw0_s1_readdata), //                    .readdata
		.in_port  (sw0_export)                         // external_connection.export
	);

	nios2e_DIP1 sw1 (
		.clk      (clk_clk),                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),   //               reset.reset_n
		.address  (mm_interconnect_0_sw1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sw1_s1_readdata), //                    .readdata
		.in_port  (sw1_export)                         // external_connection.export
	);

	nios2e_mm_interconnect_0 mm_interconnect_0 (
		.CLK_clk_clk                             (clk_clk),                                              //                           CLK_clk.clk
		.NIOS2_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                       // NIOS2_reset_reset_bridge_in_reset.reset
		.NIOS2_data_master_address               (nios2_data_master_address),                            //                 NIOS2_data_master.address
		.NIOS2_data_master_waitrequest           (nios2_data_master_waitrequest),                        //                                  .waitrequest
		.NIOS2_data_master_byteenable            (nios2_data_master_byteenable),                         //                                  .byteenable
		.NIOS2_data_master_read                  (nios2_data_master_read),                               //                                  .read
		.NIOS2_data_master_readdata              (nios2_data_master_readdata),                           //                                  .readdata
		.NIOS2_data_master_write                 (nios2_data_master_write),                              //                                  .write
		.NIOS2_data_master_writedata             (nios2_data_master_writedata),                          //                                  .writedata
		.NIOS2_data_master_debugaccess           (nios2_data_master_debugaccess),                        //                                  .debugaccess
		.NIOS2_instruction_master_address        (nios2_instruction_master_address),                     //          NIOS2_instruction_master.address
		.NIOS2_instruction_master_waitrequest    (nios2_instruction_master_waitrequest),                 //                                  .waitrequest
		.NIOS2_instruction_master_read           (nios2_instruction_master_read),                        //                                  .read
		.NIOS2_instruction_master_readdata       (nios2_instruction_master_readdata),                    //                                  .readdata
		.CYCLE_s1_address                        (mm_interconnect_0_cycle_s1_address),                   //                          CYCLE_s1.address
		.CYCLE_s1_write                          (mm_interconnect_0_cycle_s1_write),                     //                                  .write
		.CYCLE_s1_readdata                       (mm_interconnect_0_cycle_s1_readdata),                  //                                  .readdata
		.CYCLE_s1_writedata                      (mm_interconnect_0_cycle_s1_writedata),                 //                                  .writedata
		.CYCLE_s1_chipselect                     (mm_interconnect_0_cycle_s1_chipselect),                //                                  .chipselect
		.DIP0_s1_address                         (mm_interconnect_0_dip0_s1_address),                    //                           DIP0_s1.address
		.DIP0_s1_readdata                        (mm_interconnect_0_dip0_s1_readdata),                   //                                  .readdata
		.DIP1_s1_address                         (mm_interconnect_0_dip1_s1_address),                    //                           DIP1_s1.address
		.DIP1_s1_readdata                        (mm_interconnect_0_dip1_s1_readdata),                   //                                  .readdata
		.DIP2_s1_address                         (mm_interconnect_0_dip2_s1_address),                    //                           DIP2_s1.address
		.DIP2_s1_readdata                        (mm_interconnect_0_dip2_s1_readdata),                   //                                  .readdata
		.DIP3_s1_address                         (mm_interconnect_0_dip3_s1_address),                    //                           DIP3_s1.address
		.DIP3_s1_readdata                        (mm_interconnect_0_dip3_s1_readdata),                   //                                  .readdata
		.DUTY_s1_address                         (mm_interconnect_0_duty_s1_address),                    //                           DUTY_s1.address
		.DUTY_s1_write                           (mm_interconnect_0_duty_s1_write),                      //                                  .write
		.DUTY_s1_readdata                        (mm_interconnect_0_duty_s1_readdata),                   //                                  .readdata
		.DUTY_s1_writedata                       (mm_interconnect_0_duty_s1_writedata),                  //                                  .writedata
		.DUTY_s1_chipselect                      (mm_interconnect_0_duty_s1_chipselect),                 //                                  .chipselect
		.ID_control_slave_address                (mm_interconnect_0_id_control_slave_address),           //                  ID_control_slave.address
		.ID_control_slave_readdata               (mm_interconnect_0_id_control_slave_readdata),          //                                  .readdata
		.JTAG_avalon_jtag_slave_address          (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //            JTAG_avalon_jtag_slave.address
		.JTAG_avalon_jtag_slave_write            (mm_interconnect_0_jtag_avalon_jtag_slave_write),       //                                  .write
		.JTAG_avalon_jtag_slave_read             (mm_interconnect_0_jtag_avalon_jtag_slave_read),        //                                  .read
		.JTAG_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                                  .readdata
		.JTAG_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                                  .writedata
		.JTAG_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                                  .waitrequest
		.JTAG_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  //                                  .chipselect
		.LED0_s1_address                         (mm_interconnect_0_led0_s1_address),                    //                           LED0_s1.address
		.LED0_s1_write                           (mm_interconnect_0_led0_s1_write),                      //                                  .write
		.LED0_s1_readdata                        (mm_interconnect_0_led0_s1_readdata),                   //                                  .readdata
		.LED0_s1_writedata                       (mm_interconnect_0_led0_s1_writedata),                  //                                  .writedata
		.LED0_s1_chipselect                      (mm_interconnect_0_led0_s1_chipselect),                 //                                  .chipselect
		.LED1_s1_address                         (mm_interconnect_0_led1_s1_address),                    //                           LED1_s1.address
		.LED1_s1_write                           (mm_interconnect_0_led1_s1_write),                      //                                  .write
		.LED1_s1_readdata                        (mm_interconnect_0_led1_s1_readdata),                   //                                  .readdata
		.LED1_s1_writedata                       (mm_interconnect_0_led1_s1_writedata),                  //                                  .writedata
		.LED1_s1_chipselect                      (mm_interconnect_0_led1_s1_chipselect),                 //                                  .chipselect
		.LED2_s1_address                         (mm_interconnect_0_led2_s1_address),                    //                           LED2_s1.address
		.LED2_s1_write                           (mm_interconnect_0_led2_s1_write),                      //                                  .write
		.LED2_s1_readdata                        (mm_interconnect_0_led2_s1_readdata),                   //                                  .readdata
		.LED2_s1_writedata                       (mm_interconnect_0_led2_s1_writedata),                  //                                  .writedata
		.LED2_s1_chipselect                      (mm_interconnect_0_led2_s1_chipselect),                 //                                  .chipselect
		.LED3_s1_address                         (mm_interconnect_0_led3_s1_address),                    //                           LED3_s1.address
		.LED3_s1_write                           (mm_interconnect_0_led3_s1_write),                      //                                  .write
		.LED3_s1_readdata                        (mm_interconnect_0_led3_s1_readdata),                   //                                  .readdata
		.LED3_s1_writedata                       (mm_interconnect_0_led3_s1_writedata),                  //                                  .writedata
		.LED3_s1_chipselect                      (mm_interconnect_0_led3_s1_chipselect),                 //                                  .chipselect
		.LED4_s1_address                         (mm_interconnect_0_led4_s1_address),                    //                           LED4_s1.address
		.LED4_s1_write                           (mm_interconnect_0_led4_s1_write),                      //                                  .write
		.LED4_s1_readdata                        (mm_interconnect_0_led4_s1_readdata),                   //                                  .readdata
		.LED4_s1_writedata                       (mm_interconnect_0_led4_s1_writedata),                  //                                  .writedata
		.LED4_s1_chipselect                      (mm_interconnect_0_led4_s1_chipselect),                 //                                  .chipselect
		.LED5_s1_address                         (mm_interconnect_0_led5_s1_address),                    //                           LED5_s1.address
		.LED5_s1_write                           (mm_interconnect_0_led5_s1_write),                      //                                  .write
		.LED5_s1_readdata                        (mm_interconnect_0_led5_s1_readdata),                   //                                  .readdata
		.LED5_s1_writedata                       (mm_interconnect_0_led5_s1_writedata),                  //                                  .writedata
		.LED5_s1_chipselect                      (mm_interconnect_0_led5_s1_chipselect),                 //                                  .chipselect
		.LED6_s1_address                         (mm_interconnect_0_led6_s1_address),                    //                           LED6_s1.address
		.LED6_s1_write                           (mm_interconnect_0_led6_s1_write),                      //                                  .write
		.LED6_s1_readdata                        (mm_interconnect_0_led6_s1_readdata),                   //                                  .readdata
		.LED6_s1_writedata                       (mm_interconnect_0_led6_s1_writedata),                  //                                  .writedata
		.LED6_s1_chipselect                      (mm_interconnect_0_led6_s1_chipselect),                 //                                  .chipselect
		.LED7_s1_address                         (mm_interconnect_0_led7_s1_address),                    //                           LED7_s1.address
		.LED7_s1_write                           (mm_interconnect_0_led7_s1_write),                      //                                  .write
		.LED7_s1_readdata                        (mm_interconnect_0_led7_s1_readdata),                   //                                  .readdata
		.LED7_s1_writedata                       (mm_interconnect_0_led7_s1_writedata),                  //                                  .writedata
		.LED7_s1_chipselect                      (mm_interconnect_0_led7_s1_chipselect),                 //                                  .chipselect
		.NIOS2_debug_mem_slave_address           (mm_interconnect_0_nios2_debug_mem_slave_address),      //             NIOS2_debug_mem_slave.address
		.NIOS2_debug_mem_slave_write             (mm_interconnect_0_nios2_debug_mem_slave_write),        //                                  .write
		.NIOS2_debug_mem_slave_read              (mm_interconnect_0_nios2_debug_mem_slave_read),         //                                  .read
		.NIOS2_debug_mem_slave_readdata          (mm_interconnect_0_nios2_debug_mem_slave_readdata),     //                                  .readdata
		.NIOS2_debug_mem_slave_writedata         (mm_interconnect_0_nios2_debug_mem_slave_writedata),    //                                  .writedata
		.NIOS2_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_debug_mem_slave_byteenable),   //                                  .byteenable
		.NIOS2_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_debug_mem_slave_waitrequest),  //                                  .waitrequest
		.NIOS2_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_debug_mem_slave_debugaccess),  //                                  .debugaccess
		.RAM_s1_address                          (mm_interconnect_0_ram_s1_address),                     //                            RAM_s1.address
		.RAM_s1_write                            (mm_interconnect_0_ram_s1_write),                       //                                  .write
		.RAM_s1_readdata                         (mm_interconnect_0_ram_s1_readdata),                    //                                  .readdata
		.RAM_s1_writedata                        (mm_interconnect_0_ram_s1_writedata),                   //                                  .writedata
		.RAM_s1_byteenable                       (mm_interconnect_0_ram_s1_byteenable),                  //                                  .byteenable
		.RAM_s1_chipselect                       (mm_interconnect_0_ram_s1_chipselect),                  //                                  .chipselect
		.RAM_s1_clken                            (mm_interconnect_0_ram_s1_clken),                       //                                  .clken
		.SW0_s1_address                          (mm_interconnect_0_sw0_s1_address),                     //                            SW0_s1.address
		.SW0_s1_readdata                         (mm_interconnect_0_sw0_s1_readdata),                    //                                  .readdata
		.SW1_s1_address                          (mm_interconnect_0_sw1_s1_address),                     //                            SW1_s1.address
		.SW1_s1_readdata                         (mm_interconnect_0_sw1_s1_readdata)                     //                                  .readdata
	);

	nios2e_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_irq_irq)                   //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (nios2_debug_reset_request_reset),    // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
